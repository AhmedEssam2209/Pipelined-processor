LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY F_D IS
	PORT(	CLK, RST,PREV_STALL_IN: IN STD_LOGIC;
		INST: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		PC: IN STD_LOGIC_VECTOR(31 DOWNTO 0); 
		IN_PORT_IN: IN STD_LOGIC_VECTOR(31 DOWNTO 0); 
		INTERRUPT_SIG: IN STD_LOGIC;
		PREV_STALL_OUT: OUT STD_LOGIC;
		PC_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0); 
		OP_CODE: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		SRC1, SRC2, DEST: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		IN_PORT_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		INTERRUPT_SIG_OUT: OUT STD_LOGIC;
		lastpredin:in std_logic;
		lastpredOut:out std_logic





);
		
END ENTITY;

ARCHITECTURE FDREGARCH OF F_D IS
BEGIN

	PROCESS(CLK) IS
	BEGIN
	
		IF RISING_EDGE(CLK) THEN

			IF RST = '1' THEN
			OP_CODE <= (OTHERS => '0');
			PC_OUT <= (OTHERS => '0');
			SRC1 <= (OTHERS => '0');
			SRC2 <= (OTHERS => '0');
			DEST <= (OTHERS => '0');
			IN_PORT_OUT <= (OTHERS => '0');
			PREV_STALL_OUT <= '0';
			INTERRUPT_SIG_OUT <= '0';
			lastpredOut<='0';
			else
			
			OP_CODE <= INST(15 DOWNTO 11);
			SRC1 <= INST(10 DOWNTO 8); 
			SRC2 <= INST(7 DOWNTO 5);
			DEST <= INST(4 DOWNTO 2);
			lastpredOut<=lastpredin;

				
			PREV_STALL_OUT <= PREV_STALL_IN;
			IN_PORT_OUT<=IN_PORT_IN;
			INTERRUPT_SIG_OUT <= INTERRUPT_SIG;
				if INTERRUPT_SIG = '1' then
				PC_OUT <= STD_LOGIC_VECTOR(unsigned(PC) - 1 );
				else
				PC_OUT <= PC;
				end if;
			END IF; 

		END IF;
	END PROCESS;

END ARCHITECTURE;





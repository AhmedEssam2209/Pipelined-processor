LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY INSTRUCTION_CACHE IS

PORT (
CLK, RST : IN std_logic;
PC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
DATAOUT : OUT std_logic_vector(15 DOWNTO 0);
RESET_VALUE , INT_VALUE: OUT std_logic_vector(31 DOWNTO 0);
EXCEPTION_OUT : OUT STD_LOGIC 
);

END ENTITY;

ARCHITECTURE ARCH OF INSTRUCTION_CACHE IS
signal DATA : std_logic_vector(15 DOWNTO 0);
TYPE ram_type IS ARRAY(4095 DOWNTO 0) of std_logic_vector(15 DOWNTO 0);
SIGNAL INSTRUCTION_CACHE : ram_type ;

BEGIN

PROCESS(CLK) IS
BEGIN


IF FALLING_EDGE(CLK) THEN
IF to_integer(unsigned(PC))>4095 OR to_integer(unsigned(PC)) <0 THEN
EXCEPTION_OUT<= '1';
ELSE
EXCEPTION_OUT<= '0';
DATA <=INSTRUCTION_CACHE(to_integer(unsigned(PC)));
END IF;
END IF;
END PROCESS;

DATAOUT <= DATA;
RESET_VALUE <= INSTRUCTION_CACHE(1) & INSTRUCTION_CACHE(0);
INT_VALUE <= INSTRUCTION_CACHE(3) & INSTRUCTION_CACHE(2);

END ARCHITECTURE;
